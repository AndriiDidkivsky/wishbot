module parser


pub fn parse_static(options StaticParserConfig) {

}




